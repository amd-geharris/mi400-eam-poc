//=============================================================================
// AMD 2024
// All rights reserved
//
//  File Name: Top_DFX_Main.sv
//  Created By: 
//  Creation Date: September-13-2024
// 
//  Module Description:
// 
//=============================================================================    
`timescale 1 ns / 1 ns
module Top_DFX_Main #(
    //############################################################
    // Global Parameters
    //############################################################
)
(
    input AxiBusClock,
    input Clock,
    input aUART_rxd,
    output aUART_txd,
    input dReset_n,
    output [31:0]sMcuInputControl,
    input [31:0]sMcuOutputControl,
    input xAxiBusReset_n,
    input [31:0]xPcieToDfx_AXI_araddr,
    input [2:0]xPcieToDfx_AXI_arprot,
    output xPcieToDfx_AXI_arready,
    input xPcieToDfx_AXI_arvalid,
    input [31:0]xPcieToDfx_AXI_awaddr,
    input [2:0]xPcieToDfx_AXI_awprot,
    output xPcieToDfx_AXI_awready,
    input xPcieToDfx_AXI_awvalid,
    input xPcieToDfx_AXI_bready,
    output [1:0]xPcieToDfx_AXI_bresp,
    output xPcieToDfx_AXI_bvalid,
    output [31:0]xPcieToDfx_AXI_rdata,
    input xPcieToDfx_AXI_rready,
    output [1:0]xPcieToDfx_AXI_rresp,
    output xPcieToDfx_AXI_rvalid,
    input [31:0]xPcieToDfx_AXI_wdata,
    output xPcieToDfx_AXI_wready,
    input [3:0]xPcieToDfx_AXI_wstrb,
    input xPcieToDfx_AXI_wvalid
);
//=====================================================================================================================
//                                      X.X -- Local Variables
//=====================================================================================================================
//=====================================================================================================================
//                                      X.X -- Section
//=====================================================================================================================
    //############################################################
    // Micro Blaze Core
    //############################################################
    MicroBlazeCore_wrapper  MicroBlazeCore_wrapper_inst (
        .AxiBusClock(AxiBusClock),
        .Clock(Clock),
        .aUART_rxd(aUART_rxd),
        .aUART_txd(aUART_txd),
        .dReset_n(dReset_n),
        .sMcuInputControl(sMcuInputControl),
        .sMcuOutputControl(sMcuOutputControl),
        .xAxiBusReset_n(xAxiBusReset_n),
        .xPcieToDfx_AXI_araddr(xPcieToDfx_AXI_araddr),
        .xPcieToDfx_AXI_arprot(xPcieToDfx_AXI_arprot),
        .xPcieToDfx_AXI_arready(xPcieToDfx_AXI_arready),
        .xPcieToDfx_AXI_arvalid(xPcieToDfx_AXI_arvalid),
        .xPcieToDfx_AXI_awaddr(xPcieToDfx_AXI_awaddr),
        .xPcieToDfx_AXI_awprot(xPcieToDfx_AXI_awprot),
        .xPcieToDfx_AXI_awready(xPcieToDfx_AXI_awready),
        .xPcieToDfx_AXI_awvalid(xPcieToDfx_AXI_awvalid),
        .xPcieToDfx_AXI_bready(xPcieToDfx_AXI_bready),
        .xPcieToDfx_AXI_bresp(xPcieToDfx_AXI_bresp),
        .xPcieToDfx_AXI_bvalid(xPcieToDfx_AXI_bvalid),
        .xPcieToDfx_AXI_rdata(xPcieToDfx_AXI_rdata),
        .xPcieToDfx_AXI_rready(xPcieToDfx_AXI_rready),
        .xPcieToDfx_AXI_rresp(xPcieToDfx_AXI_rresp),
        .xPcieToDfx_AXI_rvalid(xPcieToDfx_AXI_rvalid),
        .xPcieToDfx_AXI_wdata(xPcieToDfx_AXI_wdata),
        .xPcieToDfx_AXI_wready(xPcieToDfx_AXI_wready),
        .xPcieToDfx_AXI_wstrb(xPcieToDfx_AXI_wstrb),
        .xPcieToDfx_AXI_wvalid(xPcieToDfx_AXI_wvalid)
    );




//=====================================================================================================================
endmodule