//=============================================================================
// AMD 2024
// All rights reserved
//
//  File Name: TopMi400EamPoc.v
//  Created By: 
//  Creation Date: August-29-2024
// 
//  Module Description:
// 
//=============================================================================
`timescale 1 ns / 1 ns

module TopMi400EamPoc
(
    // CORE
    input   wire    FPGA_CLK_100MHZ_P,
    input   wire    FPGA_CLK_100MHZ_N,
    input   wire    uMicroBlazeRst_n,

    // UART
    input   wire    MICROBLAZE_UART_RX,
    output  wire    MICROBLAZE_UART_TX

);
//=====================================================================================================================
//                                      X.X -- Local Variables
//=====================================================================================================================

//=====================================================================================================================
//                                      X.X -- Module Parameters
//=====================================================================================================================

//=====================================================================================================================
//                                      X.X -- Module Instances
//=====================================================================================================================
    //############################################################
    // Micro Blaze Core
    //############################################################
    MicroBlazeCore_wrapper MicroBlazeCore_i
        (
            .aMICROBLAZE_UART_rxd(MICROBLAZE_UART_RX),
            .aMICROBLAZE_UART_txd(MICROBLAZE_UART_TX),
            .diff_MicroBlazeClock_clk_n(FPGA_CLK_100MHZ_N),
            .diff_MicroBlazeClock_clk_p(FPGA_CLK_100MHZ_P),
            .sMcuInputControl(sMcuInputControl),
            .sMcuOutputControl(sMcuOutputControl),
            .uMicroBlazeRst_n(uMicroBlazeRst_n)
        );
//=====================================================================================================================
//                                      X.X -- Bus Assignments
//=====================================================================================================================

//=====================================================================================================================
//                                      X.X -- BiDir Assignments
//=====================================================================================================================

//=====================================================================================================================
//                                      X.X -- Input Buffers
//=====================================================================================================================

//=====================================================================================================================
//                                      X.X -- Output Assignments
//=====================================================================================================================



//=====================================================================================================================
endmodule
